magic
tech gf180mcuD
magscale 1 10
timestamp 1700892598
<< nwell >>
rect 1258 147744 238646 148262
rect 1258 146176 238646 147040
rect 1258 144608 238646 145472
rect 1258 143040 238646 143904
rect 1258 141472 238646 142336
rect 1258 139904 238646 140768
rect 1258 138336 238646 139200
rect 1258 136768 238646 137632
rect 1258 135200 238646 136064
rect 1258 133632 238646 134496
rect 1258 132064 238646 132928
rect 1258 130496 238646 131360
rect 1258 128928 238646 129792
rect 1258 127360 238646 128224
rect 1258 125792 238646 126656
rect 1258 124224 238646 125088
rect 1258 122656 238646 123520
rect 1258 121088 238646 121952
rect 1258 119545 238646 120384
rect 1258 119520 111181 119545
rect 1258 118791 121416 118816
rect 1258 117977 238646 118791
rect 1258 117952 103117 117977
rect 1258 117223 60221 117248
rect 1258 116409 238646 117223
rect 1258 116384 55853 116409
rect 1258 115655 53165 115680
rect 1258 114841 238646 115655
rect 1258 114816 32557 114841
rect 1258 114087 36589 114112
rect 1258 113273 238646 114087
rect 1258 113248 31101 113273
rect 1258 112519 30205 112544
rect 1258 111705 238646 112519
rect 1258 111680 39320 111705
rect 1258 110951 27672 110976
rect 1258 110137 238646 110951
rect 1258 110112 23709 110137
rect 1258 109383 18221 109408
rect 1258 108569 238646 109383
rect 1258 108544 17325 108569
rect 1258 107815 35719 107840
rect 1258 107001 238646 107815
rect 1258 106976 29981 107001
rect 1258 106247 26061 106272
rect 1258 105433 238646 106247
rect 1258 105408 16541 105433
rect 1258 104679 20685 104704
rect 1258 103865 238646 104679
rect 1258 103840 16429 103865
rect 1258 103111 20125 103136
rect 1258 102297 238646 103111
rect 1258 102272 25725 102297
rect 1258 101543 34573 101568
rect 1258 100729 238646 101543
rect 1258 100704 26061 100729
rect 1258 99975 19901 100000
rect 1258 99161 238646 99975
rect 1258 99136 37821 99161
rect 1258 98407 20125 98432
rect 1258 97593 238646 98407
rect 1258 97568 18333 97593
rect 1258 96839 20461 96864
rect 1258 96025 238646 96839
rect 1258 96000 18221 96025
rect 1258 95271 44541 95296
rect 1258 94457 238646 95271
rect 1258 94432 53501 94457
rect 1258 93703 14749 93728
rect 1258 92889 238646 93703
rect 1258 92864 15421 92889
rect 1258 92135 51709 92160
rect 1258 91321 238646 92135
rect 1258 91296 16317 91321
rect 1258 90567 22589 90592
rect 1258 89753 238646 90567
rect 1258 89728 15981 89753
rect 1258 88999 14637 89024
rect 1258 88185 238646 88999
rect 1258 88160 17101 88185
rect 1258 87431 33901 87456
rect 1258 86617 238646 87431
rect 1258 86592 24493 86617
rect 1258 85863 18221 85888
rect 1258 85049 238646 85863
rect 1258 85024 22477 85049
rect 1258 84295 36925 84320
rect 1258 83481 238646 84295
rect 1258 83456 23373 83481
rect 1258 82727 30093 82752
rect 1258 81913 238646 82727
rect 1258 81888 25277 81913
rect 1258 81159 20909 81184
rect 1258 80345 238646 81159
rect 1258 80320 64968 80345
rect 1258 79591 19453 79616
rect 1258 78777 238646 79591
rect 1258 78752 22141 78777
rect 1258 78023 19677 78048
rect 1258 77209 238646 78023
rect 1258 77184 26888 77209
rect 1258 76455 21917 76480
rect 1258 75641 238646 76455
rect 1258 75616 31549 75641
rect 1258 74887 21133 74912
rect 1258 74073 238646 74887
rect 1258 74048 22141 74073
rect 1258 73319 26285 73344
rect 1258 72505 238646 73319
rect 1258 72480 33944 72505
rect 1258 71751 20349 71776
rect 1258 70937 238646 71751
rect 1258 70912 22141 70937
rect 1258 70183 20349 70208
rect 1258 69369 238646 70183
rect 1258 69344 24045 69369
rect 1258 68615 28749 68640
rect 1258 67801 238646 68615
rect 1258 67776 15869 67801
rect 1258 67047 19789 67072
rect 1258 66233 238646 67047
rect 1258 66208 18445 66233
rect 1258 65479 19789 65504
rect 1258 64665 238646 65479
rect 1258 64640 31032 64665
rect 1258 63911 13853 63936
rect 1258 63097 238646 63911
rect 1258 63072 24157 63097
rect 1258 62343 14525 62368
rect 1258 61529 238646 62343
rect 1258 61504 15869 61529
rect 1258 60775 22589 60800
rect 1258 59961 238646 60775
rect 1258 59936 22141 59961
rect 1258 59207 30429 59232
rect 1258 58393 238646 59207
rect 1258 58368 18221 58393
rect 1258 57639 18221 57664
rect 1258 56825 238646 57639
rect 1258 56800 18221 56825
rect 1258 56071 12173 56096
rect 1258 55257 238646 56071
rect 1258 55232 18669 55257
rect 1258 54503 12509 54528
rect 1258 53689 238646 54503
rect 1258 53664 38941 53689
rect 1258 52935 12888 52960
rect 1258 52121 238646 52935
rect 1258 52096 45773 52121
rect 1258 51367 26061 51392
rect 1258 50553 238646 51367
rect 1258 50528 17437 50553
rect 1258 49799 18221 49824
rect 1258 48985 238646 49799
rect 1258 48960 17549 48985
rect 1258 48231 51373 48256
rect 1258 47417 238646 48231
rect 1258 47392 22141 47417
rect 1258 46663 27741 46688
rect 1258 45849 238646 46663
rect 1258 45824 26509 45849
rect 1258 45095 28301 45120
rect 1258 44281 238646 45095
rect 1258 44256 39725 44281
rect 1258 43527 49581 43552
rect 1258 42713 238646 43527
rect 1258 42688 49064 42713
rect 1258 41959 58472 41984
rect 1258 41145 238646 41959
rect 1258 41120 70749 41145
rect 1258 40391 58541 40416
rect 1258 39577 238646 40391
rect 1258 39552 57869 39577
rect 1258 38823 120141 38848
rect 1258 38009 238646 38823
rect 1258 37984 73032 38009
rect 1258 37255 75229 37280
rect 1258 36441 238646 37255
rect 1258 36416 57869 36441
rect 1258 35687 57421 35712
rect 1258 34873 238646 35687
rect 1258 34848 81389 34873
rect 1258 34119 82285 34144
rect 1258 33305 238646 34119
rect 1258 33280 92701 33305
rect 1258 32551 68328 32576
rect 1258 31737 238646 32551
rect 1258 31712 57869 31737
rect 1258 30983 68733 31008
rect 1258 30169 238646 30983
rect 1258 30144 57869 30169
rect 1258 29415 61565 29440
rect 1258 28601 238646 29415
rect 1258 28576 71197 28601
rect 1258 27847 58653 27872
rect 1258 27033 238646 27847
rect 1258 27008 57869 27033
rect 1258 26279 73101 26304
rect 1258 25465 238646 26279
rect 1258 25440 101997 25465
rect 1258 24711 82211 24736
rect 1258 23897 238646 24711
rect 1258 23872 67061 23897
rect 1258 23143 58765 23168
rect 1258 22329 238646 23143
rect 1258 22304 57869 22329
rect 1258 21575 67865 21600
rect 1258 20761 238646 21575
rect 1258 20736 102109 20761
rect 1258 20007 110181 20032
rect 1258 19193 238646 20007
rect 1258 19168 64141 19193
rect 1258 18439 60333 18464
rect 1258 17625 238646 18439
rect 1258 17600 69517 17625
rect 1258 16871 60109 16896
rect 1258 16057 238646 16871
rect 1258 16032 92701 16057
rect 1258 15303 66045 15328
rect 1258 14489 238646 15303
rect 1258 14464 63736 14489
rect 1258 13735 127981 13760
rect 1258 12921 238646 13735
rect 1258 12896 70637 12921
rect 1258 12167 88781 12192
rect 1258 11353 238646 12167
rect 1258 11328 71085 11353
rect 1258 10599 73101 10624
rect 1258 9785 238646 10599
rect 1258 9760 74600 9785
rect 1258 9031 73997 9056
rect 1258 8217 238646 9031
rect 1258 8192 87661 8217
rect 1258 7463 83405 7488
rect 1258 6649 238646 7463
rect 1258 6624 94941 6649
rect 1258 5895 100989 5920
rect 1258 5081 238646 5895
rect 1258 5056 100653 5081
rect 1258 4327 108535 4352
rect 1258 3513 238646 4327
rect 1258 3488 112973 3513
<< pwell >>
rect 1258 147040 238646 147744
rect 1258 145472 238646 146176
rect 1258 143904 238646 144608
rect 1258 142336 238646 143040
rect 1258 140768 238646 141472
rect 1258 139200 238646 139904
rect 1258 137632 238646 138336
rect 1258 136064 238646 136768
rect 1258 134496 238646 135200
rect 1258 132928 238646 133632
rect 1258 131360 238646 132064
rect 1258 129792 238646 130496
rect 1258 128224 238646 128928
rect 1258 126656 238646 127360
rect 1258 125088 238646 125792
rect 1258 123520 238646 124224
rect 1258 121952 238646 122656
rect 1258 120384 238646 121088
rect 1258 118816 238646 119520
rect 1258 117248 238646 117952
rect 1258 115680 238646 116384
rect 1258 114112 238646 114816
rect 1258 112544 238646 113248
rect 1258 110976 238646 111680
rect 1258 109408 238646 110112
rect 1258 107840 238646 108544
rect 1258 106272 238646 106976
rect 1258 104704 238646 105408
rect 1258 103136 238646 103840
rect 1258 101568 238646 102272
rect 1258 100000 238646 100704
rect 1258 98432 238646 99136
rect 1258 96864 238646 97568
rect 1258 95296 238646 96000
rect 1258 93728 238646 94432
rect 1258 92160 238646 92864
rect 1258 90592 238646 91296
rect 1258 89024 238646 89728
rect 1258 87456 238646 88160
rect 1258 85888 238646 86592
rect 1258 84320 238646 85024
rect 1258 82752 238646 83456
rect 1258 81184 238646 81888
rect 1258 79616 238646 80320
rect 1258 78048 238646 78752
rect 1258 76480 238646 77184
rect 1258 74912 238646 75616
rect 1258 73344 238646 74048
rect 1258 71776 238646 72480
rect 1258 70208 238646 70912
rect 1258 68640 238646 69344
rect 1258 67072 238646 67776
rect 1258 65504 238646 66208
rect 1258 63936 238646 64640
rect 1258 62368 238646 63072
rect 1258 60800 238646 61504
rect 1258 59232 238646 59936
rect 1258 57664 238646 58368
rect 1258 56096 238646 56800
rect 1258 54528 238646 55232
rect 1258 52960 238646 53664
rect 1258 51392 238646 52096
rect 1258 49824 238646 50528
rect 1258 48256 238646 48960
rect 1258 46688 238646 47392
rect 1258 45120 238646 45824
rect 1258 43552 238646 44256
rect 1258 41984 238646 42688
rect 1258 40416 238646 41120
rect 1258 38848 238646 39552
rect 1258 37280 238646 37984
rect 1258 35712 238646 36416
rect 1258 34144 238646 34848
rect 1258 32576 238646 33280
rect 1258 31008 238646 31712
rect 1258 29440 238646 30144
rect 1258 27872 238646 28576
rect 1258 26304 238646 27008
rect 1258 24736 238646 25440
rect 1258 23168 238646 23872
rect 1258 21600 238646 22304
rect 1258 20032 238646 20736
rect 1258 18464 238646 19168
rect 1258 16896 238646 17600
rect 1258 15328 238646 16032
rect 1258 13760 238646 14464
rect 1258 12192 238646 12896
rect 1258 10624 238646 11328
rect 1258 9056 238646 9760
rect 1258 7488 238646 8192
rect 1258 5920 238646 6624
rect 1258 4352 238646 5056
rect 1258 3050 238646 3488
<< obsm1 >>
rect 1344 3076 238560 148236
<< metal2 >>
rect 6944 0 7056 800
rect 10080 0 10192 800
rect 13216 0 13328 800
rect 16352 0 16464 800
rect 19488 0 19600 800
rect 22624 0 22736 800
rect 25760 0 25872 800
rect 28896 0 29008 800
rect 32032 0 32144 800
rect 35168 0 35280 800
rect 38304 0 38416 800
rect 41440 0 41552 800
rect 44576 0 44688 800
rect 47712 0 47824 800
rect 50848 0 50960 800
rect 53984 0 54096 800
rect 57120 0 57232 800
rect 60256 0 60368 800
rect 63392 0 63504 800
rect 66528 0 66640 800
rect 69664 0 69776 800
rect 72800 0 72912 800
rect 75936 0 76048 800
rect 79072 0 79184 800
rect 82208 0 82320 800
rect 85344 0 85456 800
rect 88480 0 88592 800
rect 91616 0 91728 800
rect 94752 0 94864 800
rect 97888 0 98000 800
rect 101024 0 101136 800
rect 104160 0 104272 800
rect 107296 0 107408 800
rect 110432 0 110544 800
rect 113568 0 113680 800
rect 116704 0 116816 800
rect 119840 0 119952 800
rect 122976 0 123088 800
rect 126112 0 126224 800
rect 129248 0 129360 800
rect 132384 0 132496 800
rect 135520 0 135632 800
rect 138656 0 138768 800
rect 141792 0 141904 800
rect 144928 0 145040 800
rect 148064 0 148176 800
rect 151200 0 151312 800
rect 154336 0 154448 800
rect 157472 0 157584 800
rect 160608 0 160720 800
rect 163744 0 163856 800
rect 166880 0 166992 800
rect 170016 0 170128 800
rect 173152 0 173264 800
rect 176288 0 176400 800
rect 179424 0 179536 800
rect 182560 0 182672 800
rect 185696 0 185808 800
rect 188832 0 188944 800
rect 191968 0 192080 800
rect 195104 0 195216 800
rect 198240 0 198352 800
rect 201376 0 201488 800
rect 204512 0 204624 800
rect 207648 0 207760 800
rect 210784 0 210896 800
rect 213920 0 214032 800
rect 217056 0 217168 800
rect 220192 0 220304 800
rect 223328 0 223440 800
rect 226464 0 226576 800
rect 229600 0 229712 800
rect 232736 0 232848 800
<< obsm2 >>
rect 4476 860 236292 148214
rect 4476 130 6884 860
rect 7116 130 10020 860
rect 10252 130 13156 860
rect 13388 130 16292 860
rect 16524 130 19428 860
rect 19660 130 22564 860
rect 22796 130 25700 860
rect 25932 130 28836 860
rect 29068 130 31972 860
rect 32204 130 35108 860
rect 35340 130 38244 860
rect 38476 130 41380 860
rect 41612 130 44516 860
rect 44748 130 47652 860
rect 47884 130 50788 860
rect 51020 130 53924 860
rect 54156 130 57060 860
rect 57292 130 60196 860
rect 60428 130 63332 860
rect 63564 130 66468 860
rect 66700 130 69604 860
rect 69836 130 72740 860
rect 72972 130 75876 860
rect 76108 130 79012 860
rect 79244 130 82148 860
rect 82380 130 85284 860
rect 85516 130 88420 860
rect 88652 130 91556 860
rect 91788 130 94692 860
rect 94924 130 97828 860
rect 98060 130 100964 860
rect 101196 130 104100 860
rect 104332 130 107236 860
rect 107468 130 110372 860
rect 110604 130 113508 860
rect 113740 130 116644 860
rect 116876 130 119780 860
rect 120012 130 122916 860
rect 123148 130 126052 860
rect 126284 130 129188 860
rect 129420 130 132324 860
rect 132556 130 135460 860
rect 135692 130 138596 860
rect 138828 130 141732 860
rect 141964 130 144868 860
rect 145100 130 148004 860
rect 148236 130 151140 860
rect 151372 130 154276 860
rect 154508 130 157412 860
rect 157644 130 160548 860
rect 160780 130 163684 860
rect 163916 130 166820 860
rect 167052 130 169956 860
rect 170188 130 173092 860
rect 173324 130 176228 860
rect 176460 130 179364 860
rect 179596 130 182500 860
rect 182732 130 185636 860
rect 185868 130 188772 860
rect 189004 130 191908 860
rect 192140 130 195044 860
rect 195276 130 198180 860
rect 198412 130 201316 860
rect 201548 130 204452 860
rect 204684 130 207588 860
rect 207820 130 210724 860
rect 210956 130 213860 860
rect 214092 130 216996 860
rect 217228 130 220132 860
rect 220364 130 223268 860
rect 223500 130 226404 860
rect 226636 130 229540 860
rect 229772 130 232676 860
rect 232908 130 236292 860
<< obsm3 >>
rect 4466 28 235150 148204
<< metal4 >>
rect 4448 3076 4768 148236
rect 19808 3076 20128 148236
rect 35168 3076 35488 148236
rect 50528 3076 50848 148236
rect 65888 3076 66208 148236
rect 81248 3076 81568 148236
rect 96608 3076 96928 148236
rect 111968 3076 112288 148236
rect 127328 3076 127648 148236
rect 142688 3076 143008 148236
rect 158048 3076 158368 148236
rect 173408 3076 173728 148236
rect 188768 3076 189088 148236
rect 204128 3076 204448 148236
rect 219488 3076 219808 148236
rect 234848 3076 235168 148236
<< obsm4 >>
rect 20748 3016 35108 129678
rect 35548 3016 50468 129678
rect 50908 3016 65828 129678
rect 66268 3016 81188 129678
rect 81628 3016 96548 129678
rect 96988 3016 111908 129678
rect 112348 3016 127268 129678
rect 127708 3016 142628 129678
rect 143068 3016 157988 129678
rect 158428 3016 173348 129678
rect 173788 3016 188708 129678
rect 189148 3016 204068 129678
rect 204508 3016 205044 129678
rect 20748 18 205044 3016
<< labels >>
rlabel metal2 s 13216 0 13328 800 6 la_data_in[0]
port 1 nsew signal input
rlabel metal2 s 75936 0 76048 800 6 la_data_in[10]
port 2 nsew signal input
rlabel metal2 s 82208 0 82320 800 6 la_data_in[11]
port 3 nsew signal input
rlabel metal2 s 88480 0 88592 800 6 la_data_in[12]
port 4 nsew signal input
rlabel metal2 s 94752 0 94864 800 6 la_data_in[13]
port 5 nsew signal input
rlabel metal2 s 101024 0 101136 800 6 la_data_in[14]
port 6 nsew signal input
rlabel metal2 s 107296 0 107408 800 6 la_data_in[15]
port 7 nsew signal input
rlabel metal2 s 113568 0 113680 800 6 la_data_in[16]
port 8 nsew signal input
rlabel metal2 s 119840 0 119952 800 6 la_data_in[17]
port 9 nsew signal input
rlabel metal2 s 126112 0 126224 800 6 la_data_in[18]
port 10 nsew signal input
rlabel metal2 s 132384 0 132496 800 6 la_data_in[19]
port 11 nsew signal input
rlabel metal2 s 19488 0 19600 800 6 la_data_in[1]
port 12 nsew signal input
rlabel metal2 s 138656 0 138768 800 6 la_data_in[20]
port 13 nsew signal input
rlabel metal2 s 144928 0 145040 800 6 la_data_in[21]
port 14 nsew signal input
rlabel metal2 s 151200 0 151312 800 6 la_data_in[22]
port 15 nsew signal input
rlabel metal2 s 157472 0 157584 800 6 la_data_in[23]
port 16 nsew signal input
rlabel metal2 s 163744 0 163856 800 6 la_data_in[24]
port 17 nsew signal input
rlabel metal2 s 170016 0 170128 800 6 la_data_in[25]
port 18 nsew signal input
rlabel metal2 s 176288 0 176400 800 6 la_data_in[26]
port 19 nsew signal input
rlabel metal2 s 182560 0 182672 800 6 la_data_in[27]
port 20 nsew signal input
rlabel metal2 s 188832 0 188944 800 6 la_data_in[28]
port 21 nsew signal input
rlabel metal2 s 195104 0 195216 800 6 la_data_in[29]
port 22 nsew signal input
rlabel metal2 s 25760 0 25872 800 6 la_data_in[2]
port 23 nsew signal input
rlabel metal2 s 201376 0 201488 800 6 la_data_in[30]
port 24 nsew signal input
rlabel metal2 s 207648 0 207760 800 6 la_data_in[31]
port 25 nsew signal input
rlabel metal2 s 213920 0 214032 800 6 la_data_in[32]
port 26 nsew signal input
rlabel metal2 s 217056 0 217168 800 6 la_data_in[33]
port 27 nsew signal input
rlabel metal2 s 220192 0 220304 800 6 la_data_in[34]
port 28 nsew signal input
rlabel metal2 s 223328 0 223440 800 6 la_data_in[35]
port 29 nsew signal input
rlabel metal2 s 226464 0 226576 800 6 la_data_in[36]
port 30 nsew signal input
rlabel metal2 s 229600 0 229712 800 6 la_data_in[37]
port 31 nsew signal input
rlabel metal2 s 232736 0 232848 800 6 la_data_in[38]
port 32 nsew signal input
rlabel metal2 s 32032 0 32144 800 6 la_data_in[3]
port 33 nsew signal input
rlabel metal2 s 38304 0 38416 800 6 la_data_in[4]
port 34 nsew signal input
rlabel metal2 s 44576 0 44688 800 6 la_data_in[5]
port 35 nsew signal input
rlabel metal2 s 50848 0 50960 800 6 la_data_in[6]
port 36 nsew signal input
rlabel metal2 s 57120 0 57232 800 6 la_data_in[7]
port 37 nsew signal input
rlabel metal2 s 63392 0 63504 800 6 la_data_in[8]
port 38 nsew signal input
rlabel metal2 s 69664 0 69776 800 6 la_data_in[9]
port 39 nsew signal input
rlabel metal2 s 16352 0 16464 800 6 la_data_out[0]
port 40 nsew signal output
rlabel metal2 s 79072 0 79184 800 6 la_data_out[10]
port 41 nsew signal output
rlabel metal2 s 85344 0 85456 800 6 la_data_out[11]
port 42 nsew signal output
rlabel metal2 s 91616 0 91728 800 6 la_data_out[12]
port 43 nsew signal output
rlabel metal2 s 97888 0 98000 800 6 la_data_out[13]
port 44 nsew signal output
rlabel metal2 s 104160 0 104272 800 6 la_data_out[14]
port 45 nsew signal output
rlabel metal2 s 110432 0 110544 800 6 la_data_out[15]
port 46 nsew signal output
rlabel metal2 s 116704 0 116816 800 6 la_data_out[16]
port 47 nsew signal output
rlabel metal2 s 122976 0 123088 800 6 la_data_out[17]
port 48 nsew signal output
rlabel metal2 s 129248 0 129360 800 6 la_data_out[18]
port 49 nsew signal output
rlabel metal2 s 135520 0 135632 800 6 la_data_out[19]
port 50 nsew signal output
rlabel metal2 s 22624 0 22736 800 6 la_data_out[1]
port 51 nsew signal output
rlabel metal2 s 141792 0 141904 800 6 la_data_out[20]
port 52 nsew signal output
rlabel metal2 s 148064 0 148176 800 6 la_data_out[21]
port 53 nsew signal output
rlabel metal2 s 154336 0 154448 800 6 la_data_out[22]
port 54 nsew signal output
rlabel metal2 s 160608 0 160720 800 6 la_data_out[23]
port 55 nsew signal output
rlabel metal2 s 166880 0 166992 800 6 la_data_out[24]
port 56 nsew signal output
rlabel metal2 s 173152 0 173264 800 6 la_data_out[25]
port 57 nsew signal output
rlabel metal2 s 179424 0 179536 800 6 la_data_out[26]
port 58 nsew signal output
rlabel metal2 s 185696 0 185808 800 6 la_data_out[27]
port 59 nsew signal output
rlabel metal2 s 191968 0 192080 800 6 la_data_out[28]
port 60 nsew signal output
rlabel metal2 s 198240 0 198352 800 6 la_data_out[29]
port 61 nsew signal output
rlabel metal2 s 28896 0 29008 800 6 la_data_out[2]
port 62 nsew signal output
rlabel metal2 s 204512 0 204624 800 6 la_data_out[30]
port 63 nsew signal output
rlabel metal2 s 210784 0 210896 800 6 la_data_out[31]
port 64 nsew signal output
rlabel metal2 s 35168 0 35280 800 6 la_data_out[3]
port 65 nsew signal output
rlabel metal2 s 41440 0 41552 800 6 la_data_out[4]
port 66 nsew signal output
rlabel metal2 s 47712 0 47824 800 6 la_data_out[5]
port 67 nsew signal output
rlabel metal2 s 53984 0 54096 800 6 la_data_out[6]
port 68 nsew signal output
rlabel metal2 s 60256 0 60368 800 6 la_data_out[7]
port 69 nsew signal output
rlabel metal2 s 66528 0 66640 800 6 la_data_out[8]
port 70 nsew signal output
rlabel metal2 s 72800 0 72912 800 6 la_data_out[9]
port 71 nsew signal output
rlabel metal4 s 4448 3076 4768 148236 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 148236 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 148236 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 148236 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 148236 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 148236 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 148236 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 219488 3076 219808 148236 6 vdd
port 72 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 148236 6 vss
port 73 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 148236 6 vss
port 73 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 148236 6 vss
port 73 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 148236 6 vss
port 73 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 148236 6 vss
port 73 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 148236 6 vss
port 73 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 148236 6 vss
port 73 nsew ground bidirectional
rlabel metal4 s 234848 3076 235168 148236 6 vss
port 73 nsew ground bidirectional
rlabel metal2 s 6944 0 7056 800 6 wb_clk_i
port 74 nsew signal input
rlabel metal2 s 10080 0 10192 800 6 wb_rst_i
port 75 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 240000 152000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17191366
string GDS_FILE /home/axios/Workspaces/caravel_gfmpw-1/GFMPW-1_test/openlane/present_gf180_wrapper/runs/23_11_25_13_01/results/signoff/present_gf180_wrapper.magic.gds
string GDS_START 384900
<< end >>

